
module Pipeline_CPU( clk_i, rst_n );
		
//I/O port
input         clk_i;
input         rst_n;

//Internal Signles
wire [16-1:0] PC_in;            //
wire [16-1:0] PC_ReadAddress;   //
wire [16-1:0] PCadder1_sum;     //
wire [16-1:0] PCadder2_sum;
wire [16-1:0] Instruction;      //
wire  [3-1:0] RDaddr;
wire [16-1:0] RDdata;
wire [16-1:0] RSdata;
wire [16-1:0] RTdata;

//Decoder
wire 	        RegDst;
wire 		RegWrite;
wire	[2-1:0] ALUOp;
wire	        ALUSrc;
wire	        Branch;
wire		MemtoReg;
wire		BranchType;
wire		Jump;
wire		MemRead;
wire		MemWrite;

//AC
wire  [4-1:0] ALU_operation;
wire  [2-1:0] FUResult_Select;
wire [16-1:0] FUResult;

//ALU
wire [16-1:0] SignExtend; 
wire [16-1:0] ALU_src2;
wire Zero;
wire _Zero;
wire Overflow;
wire [16-1:0] ALU_result;

//DM
wire [16-1:0] Mem_Readdata;

//branch
wire ZERO;

wire PCSrc;

//ZF
wire [16-1:0] Zerofilled;

//shifter
wire [16-1:0] Shifter_result;

//PC
wire [16-1:0] SE_shiftleft1;
wire [16-1:0] PC_branch;
wire [16-1:0] PC_jump;


//IF_ID
wire [15:0] IF_ID_Instruction;
wire [15:0] IF_ID_PCadder1_sum;

//ID_EX
wire [6:0]  ID_EX_EX ;
wire [1:0]  ID_EX_MEM ; 
wire [1:0]  ID_EX_WB ;
wire [12:0]  ID_EX_Jump_dst ; 
wire [15:0]  ID_EX_PCadder1_sum ; 
wire [15:0]  ID_EX_RSdata ;
wire [15:0]  ID_EX_RTdata ; 
wire [15:0]  ID_EX_SignExtend ; 
wire [15:0]  ID_EX_Zerofilled ; 
wire [3:0]  ID_EX_Func ;
wire [2:0]  ID_EX_RT_reg ; 
wire [2:0]  ID_EX_RD_reg ;
wire [2:0]  ID_EX_RS_reg;

wire [2:0]   Forward_A ;
wire [2:0]   Forward_B ;
wire [15:0]  Forward_A_out;
wire [15:0]  Forward_B_out;

//EX_MEM
wire [1:0] EX_MEM_WB ;
wire [1:0] EX_MEM_MEM ; 
wire [15:0] EX_MEM_FUResult ;
wire [15:0] EX_MEM_RTdata ;
wire [2:0] EX_MEM_RDaddr;
wire [2:0] EX_MEM_RTaddr;
wire      Mem_Forward;

//MEM_WB
wire [1:0] MEM_WB_WB ;
wire [15:0] MEM_WB_Mem_Readdata ;
wire [15:0] MEM_WB_FUResult;
wire [2:0] MEM_WB_RDaddr;
wire [15:0] MEM_Forward_out ;

//data_hazard_detecor
wire [15:0] PC_Const;
wire IF_ID_Hold ;
wire IF_ID_Flush;
wire Data_ID_EX_Flush;
wire PC_Hold;

// Branch_Detector
wire  Branch_ID_EX_Flush;


//module

/////////////////////////////////////////////////////////////////////////////////////////////////////////// Branch
Mux2to1 branch( PCadder1_sum ,                             ///
                PCadder2_sum ,                             ///
                PCSrc ,                                    ///
                PC_branch);                                ///
//////////////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////////////////////////////// Jump
Mux2to1 jump( PC_branch ,                                  ///
              PC_jump ,                                    ///
              ID_EX_EX[0] ,                                ///
              PC_in);                                      ///
//////////////////////////////////////////////////////////////////////////////////////////////////////////


//////////////////////////////////////////////////////////////////////////////////////////////////////////// PC
Program_Counter PC(                                        ///
        .clk_i(clk_i),                                     ///
        .rst_n(rst_n),                                     ///
        .pc_in_i(PC_in) ,                                  ///
        .pc_out_o(PC_ReadAddress)                          ///
        );                                                 ///
///////////////////////////////////////////////////////////////////////////////////////////////////////////


//////////////////////////////////////////////////////////////////////////////////////////////////////////  PCadder_1
Adder PCadder1( PC_ReadAddress ,                           /// 
                PC_Const ,                                 ///
                PCadder1_sum);                             ///
/////////////////////////////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////////////////////////  PC_Const
Mux2to1 pc_const( 16'b0000_0000_0000_0010 ,           ///
                  16'b0000_0000_0000_0000 ,           ///
                  PC_Hold ,                              ///
                  PC_Const);                             ///
 //////////////////////////////////////////////////////////////////////////////////////////////////////                

//////////////////////////////////////////////////////////////////////////////////////////////////// IM	
Instr_Memory IM(                                       ///
        .pc_addr_i(PC_ReadAddress),                    ///
        .instr_o(Instruction)                          ///
        );                                             ///
///////////////////////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////////////////////     IF_ID_Stage   ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
IF_ID_Stage IF_ID( clk_i, 
                   rst_n , 
                 
                   PCadder1_sum , 
                   Instruction , 
                   IF_ID_Hold , 
                   IF_ID_Flush ,
                   
                   IF_ID_PCadder1_sum , 
                   IF_ID_Instruction) ;
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////  Load_Use_Hazard
Load_Use_HazardDetector load_use_hazard(                                       ///
                                 .MemWrite(MemWrite) ,                         ///
                                 .ID_EX_MemRead(ID_EX_MEM[0]) ,                ///
                                 .RDaddr(RDaddr ),                             ///
                                 .IF_ID_RS(IF_ID_Instruction[12:10]) ,         ///
                                 .IF_ID_RT(IF_ID_Instruction[9:7]) ,           ///
                                 .PC_Hold(PC_Hold) ,                           ///
                                 .IF_ID_Hold(IF_ID_Hold ),                     ///
                                 .ID_EX_Flush(Data_ID_EX_Flush)) ;             ///
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////



//////////////////////////////////////////////////////////////////////////////////////// Regster
Reg_File RF(                                    ///
        .clk_i(clk_i),                          ///
	    .rst_n(rst_n) ,                         ///
        .RSaddr_i(IF_ID_Instruction[12:10]) ,   ///
        .RTaddr_i(IF_ID_Instruction[9:7]) ,     ///
        .RDaddr_i(MEM_WB_RDaddr) ,              ///
        .RDdata_i(RDdata)  ,                    ///
        .RegWrite_i(MEM_WB_WB[0]),              ///
        .RSdata_o(RSdata) ,                     ///
        .RTdata_o(RTdata)                       ///
        );                                      ///
//////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////// Decoder
Decoder decoder( IF_ID_Instruction[15:13],     ///
                 RegWrite,	                   ///
                 ALUOp,                        ///
                 ALUSrc,                       ///
                 RegDst,                       ///
                 Branch,                       ///
                 BranchType,                   ///
                 MemToReg,                     ///
                 MemRead,                      ///
                 MemWrite,                     ///
                 Jump ) ;                      ///
                                               ///
//////////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////////////////// SignExtend
Sign_Extend sign_extend( IF_ID_Instruction[6:0] ,    ///
                         SignExtend) ;               ///
/////////////////////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////////////////// Zerofilled
Zero_Filled zero_filled( IF_ID_Instruction[6:0] ,    ///
                         Zerofilled );               ///
/////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////////////////////////////     ID_EX_Stage    //////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
ID_EX_Stage  ID_EX( .clk_i(clk_i) , 
                    .rst_n(rst_n) , 
                    
                    .Data_ID_EX_Flush(Data_ID_EX_Flush) , 
                    .Branch_ID_EX_Flush(Branch_ID_EX_Flush ) ,
                    
                    .EX({ RegDst , ALUOp , ALUSrc , BranchType , Branch , Jump} ),  //EX
                    .MEM({ MemWrite , MemRead}) ,                                    //MEM
                    .WB({ MemToReg , RegWrite} ),                                   //WB
                    .jump_dst(IF_ID_Instruction[12:0]) ,
                    .PC(IF_ID_PCadder1_sum ), 
                    .RS_data(RSdata) , 
                    .RT_data(RTdata) , 
                    .SE(SignExtend) , 
                    .Zerofilled(Zerofilled) ,  
                    .func(IF_ID_Instruction[3:0]) ,
                    .RS_reg(IF_ID_Instruction[12:10] ), 
                    .RT_reg(IF_ID_Instruction[9:7]) ,
                    .RD_reg(IF_ID_Instruction[6:4]),
                    
                    .EX_o(ID_EX_EX) , 
                    .MEM_o(ID_EX_MEM) , 
                    .WB_o(ID_EX_WB) ,
                    .jump_dst_o(ID_EX_Jump_dst), 
                    .PC_o(ID_EX_PCadder1_sum) , 
                    .RS_data_o(ID_EX_RSdata) , 
                    .RT_data_o(ID_EX_RTdata) , 
                    .SE_o(ID_EX_SignExtend) , 
                    .Zerofilled_o(ID_EX_Zerofilled), 
                    .func_o(ID_EX_Func) ,
                    .RT_reg_o(ID_EX_RT_reg) , 
                    .RD_reg_o(ID_EX_RD_reg) ,
                    .RS_reg_o(ID_EX_RS_reg) );
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////////////  Data_Forwarding
EX_ForwardingUnit EX_Forwarding( EX_MEM_RDaddr , ///
                              MEM_WB_RDaddr ,    ///
                              ID_EX_RS_reg ,     ///
                              ID_EX_RT_reg ,     ///
                              EX_MEM_WB[0] ,     ///
                              MEM_WB_WB[0] ,     ///
                              Forward_A ,        ///
                              Forward_B );       ///
/////////////////////////////////////////////////////////////////////////////////////////


//////////////////////////////////////////////////////////////////////////////////////////////////////// Branch_detector
Control_Hazard_Detector control_hazard_detector( PCSrc ,  ///
                                 ID_EX_EX[0] ,            ///
                                 IF_ID_Flush ,            ///
                                 Branch_ID_EX_Flush);     ///
////////////////////////////////////////////////////////////////////////////////////////////////////////


////////////////////////////////////////////////////////////////////////////////////////// RegDst
Mux2to1_3bits Regdst( ID_EX_RT_reg ,             ///
                      ID_EX_RD_reg ,             ///
                      ID_EX_EX[6] ,              ///
                      RDaddr);                   ///
///////////////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////////////// Forward_A
Mux3to1 forward_A(  ID_EX_RSdata ,                ///  0 RS
                     RDdata ,                     ///  1 from MEM
                     EX_MEM_FUResult ,            ///  2 from EX
                    Forward_A ,                   ///
                     Forward_A_out );             ///
//////////////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////////////// Forward_B
Mux3to1 forward_B(  ID_EX_RTdata ,                ///  0  RT
                     RDdata ,                     ///  1  from MEM
                     EX_MEM_FUResult ,            ///  2  from  EX
                    Forward_B,                    ///
                    Forward_B_out  );             ///
//////////////////////////////////////////////////////////////////////////////////////////


/////////////////////////////////////////////////////////////////////////////////////////// ALU_Src
Mux2to1 ALU_Src( Forward_B_out,                   ///
                 ID_EX_SignExtend ,               ///
                 ID_EX_EX[3] ,                    ///
                 ALU_src2);                       ///
//////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////////// ALU_Ctrl
ALU_Ctrl ALU_ctrl( ID_EX_Func,                 ///
                   ID_EX_EX[5:4],              ///
                   ALU_operation,              ///
                   FUResult_Select );          ///
/////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////////////////////////////////// Shift_left_one
Shift_Left_one shift_left_one( ID_EX_SignExtend ,            ///
                  SE_shiftleft1);                            ///
//////////////////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////////// PCadder_2
Adder PCadder_2( ID_EX_PCadder1_sum ,          ///
                 SE_shiftleft1 ,               ///
                 PCadder2_sum);                ///
//////////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////// ALU
ALU alu( Forward_A_out,                        ///
         ALU_src2 ,                           ///
         ALU_operation ,                      ///
         ALU_result ,                         ///
         Zero ,                               ///
         Overflow);                           ///
////////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////// Shifter
Shifter shifter( Shifter_result ,             ///
                 ALU_operation[0] ,           ///
                 ALU_src2);                   ///
///////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////// BranchType
assign _Zero = ~Zero;                        ///
Mux2to1_1bit Branchtype( Zero ,             ///
                         _Zero ,            ///
                         ID_EX_EX[2] ,      ///
                         ZERO);             ///
/////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////// FUresult
Mux3to1 Furesult( ALU_result ,              ///
                  Shifter_result ,          ///
                  ID_EX_Zerofilled ,        ///
                  FUResult_Select ,         ///
                  FUResult);                ///
////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////// Branch_and
assign PCSrc = ZERO & ID_EX_EX[1];         ///
//////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////// Jump_assemble
assign PC_jump = { ID_EX_PCadder1_sum[15:14] , ID_EX_Jump_dst , 1'b0};     ///
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////



////////////////////////////////////////////////////////////////////////////////////////////////////////////   EX_MEM_Stage   ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
EX_MEM_Stage EX_MEM( .clk_i(clk_i) , 
                     .rst_n(rst_n) , 
                     
                     .WB(ID_EX_WB) , 
                     .MEM(ID_EX_MEM) , 
                     .FU_result(FUResult) , 
                     .RT_data(Forward_B_out) , 
                     .Write_dst(RDaddr) , 
                     .RT_addr(ID_EX_RT_reg) ,
                                      
                     .WB_o(EX_MEM_WB) , 
                     .MEM_o(EX_MEM_MEM) , 
                     .FU_result_o(EX_MEM_FUResult) , 
                     .RT_data_o(EX_MEM_RTdata), 
                     .Write_dst_o(EX_MEM_RDaddr) ,
                     .RT_addr_o(EX_MEM_RTaddr));
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////  Load_Store_Forwarding
MEM_ForwardingUnit MEM_Forwarding( MEM_WB_WB[1] ,                ///
                                          EX_MEM_MEM[1] ,        ///
                                          EX_MEM_RTaddr ,        ///
                                          MEM_WB_RDaddr ,        ///
                                          MEM_Forward );         ///
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////// MEM_Forward
Mux2to1 mem_forward( EX_MEM_RTdata ,          ///
                     RDdata ,                 ///
                     MEM_Forward ,            ///
                     MEM_Forward_out);        ///
////////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////////////////////////// Mem
Data_Memory DM(                                           ///
        .clk_i(clk_i),                                    ///
        .addr_i(EX_MEM_FUResult),                         ///
        .data_i(MEM_Forward_out),                         ///
        .MemRead_i(EX_MEM_MEM[0]),                        ///
        .MemWrite_i(EX_MEM_MEM[1]),                       ///
        .data_o(Mem_Readdata)                             ///
        );                                                ///
/////////////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////////////////////////////////////  MEM_WB_Stage /////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
MEM_WB_Stage MEM_WB( clk_i , 
                     rst_n ,
                     
                     EX_MEM_WB , 
                     Mem_Readdata , 
                     EX_MEM_FUResult , 
                     EX_MEM_RDaddr ,
                                       
                     MEM_WB_WB , 
                     MEM_WB_Mem_Readdata , 
                     MEM_WB_FUResult,
                     MEM_WB_RDaddr);
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////// MemtoReg
Mux2to1 memtoreg( MEM_WB_FUResult ,        ///
                  MEM_WB_Mem_Readdata ,    ///
                  MEM_WB_WB[1] ,           ///
                  RDdata);                 ///
///////////////////////////////////////////////////////////////////////////////             


                
 
 

endmodule

